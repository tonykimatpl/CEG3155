LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY eightBitShiftRegisterRight IS
	PORT(
		i_resetBar, i_load: STD_LOGIC;
		i_clk: IN STD_LOGIC;
		i_Value: IN STD_LOGIC_VECTOR(7 downto 0);
		o_Value: OUT STD_LOGIC_VECTOR(7 downto 0));
END eightBitShiftRegisterRight;
	
ARCHITECTURE behavior OF eightBitShiftRegisterRight IS
	SIGNAL int_Value, int_notValue: STD_LOGIC_VECTOR(7 downto 0);
	
	COMPONENT enRdFF_2
		PORT(
			i_resetBar: IN STD_LOGIC;
			i_d: IN STD_LOGIC;
			i_enable: IN STD_LOGIC;
			i_clk: IN STD_LOGIC;
			o_q, o_qBar: OUT STD_LOGIC);
	END COMPONENT;
	
BEGIN

msb:enRdFF_2
	PORT MAP (i_resetBar => i_resetBar,
	i_d => i_Value(0),
	i_enable => i_load,
	i_clk => i_clk,
	o_q => int_Value(7),
	o_qBar => int_notValue(7));
	
ssb6:enRdFF_2
	PORT MAP (i_resetBar => i_resetBar,
	i_d => int_Value(7),
	i_enable => i_load,
	i_clk => i_clk,
	o_q => int_Value(6),
	o_qBar => int_notValue(6));
	
ssb5:enRdFF_2
	PORT MAP (i_resetBar => i_resetBar,
	i_d => int_Value(6),
	i_enable => i_load,
	i_clk => i_clk,
	o_q => int_Value(5),
	o_qBar => int_notValue(5));
	
ssb4:enRdFF_2
	PORT MAP (i_resetBar => i_resetBar,
	i_d => int_Value(5),
	i_enable => i_load,
	i_clk => i_clk,
	o_q => int_Value(4),
	o_qBar => int_notValue(4));
	
ssb3:enRdFF_2
	PORT MAP (i_resetBar => i_resetBar,
	i_d => int_Value(4),
	i_enable => i_load,
	i_clk => i_clk,
	o_q => int_Value(3),
	o_qBar => int_notValue(3));
	
ssb2:enRdFF_2
	PORT MAP (i_resetBar => i_resetBar,
	i_d => int_Value(3),
	i_enable => i_load,
	i_clk => i_clk,
	o_q => int_Value(2),
	o_qBar => int_notValue(2));
	
ssb1:enRdFF_2
	PORT MAP (i_resetBar => i_resetBar,
	i_d => int_Value(2),
	i_enable => i_load,
	i_clk => i_clk,
	o_q => int_Value(1),
	o_qBar => int_notValue(1));
	
lsb:enRdFF_2
	PORT MAP (i_resetBar => i_resetBar,
	i_d => int_Value(1),
	i_enable => i_load,
	i_clk => i_clk,
	o_q => int_Value(0),
	o_qBar => int_notValue(0));
	
-- Output Driver
	o_Value		<= int_Value;

END behavior;
	
	
	
	
	
	